// Outputs a 1 for a single clock cycle when a button is pushed, "cleaning" the button input

// Copyright (C) 2023  OmarElfouly, iRustom, BavlyRemon, omaranwar1

// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.

// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.

// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.


module pushButtonDetector( clk, rst, uncleanInput, cleanOutput);
    input wire clk;
    input wire rst;
    input wire uncleanInput;
    output wire cleanOutput;

    wire newclk;
    clockDivider #(5000) newclkDiv(.clk(clk),.rst(rst) ,.clk_out(newclk));
    
    wire postBounce; 
    debouncer d(.clk(newclk),.rst(rst),.in(uncleanInput),.out(postBounce));
    
    wire postSynch;
    synchronizer s(.clk(newclk),.sig(postBounce),.sig1(postSynch));
    
    risingEdgeDetector r(.clk(newclk), .level(postSynch),.tick(cleanOutput));
    
endmodule 